***************************************
*** GAGABIRO VALVE POWER AMPLIFIER 	***
***	AUTHOR:  JOAO CARLET			***
*** CONTACT: JVCCARLET@USP.BR		***
***************************************

*RESISTORS
R1 		0 		N023 	{int(X1)*1R}
R2 		N021 	V_PP 	{int(X2)*1R}
R3 		0 		N010 	{int(X3)*1R}
R4 		N008 	V_PP 	{int(X4)*1R}
R5 		N003 	V_PP 	{int(X5)*1R}
R6 		N009 	N017 	{int(X6)*1R}
R7 		V_in 	N017 	{int(X7)*1R}
R8 		N010 	N011 	{int(X8)*1R}
R9 		0 		N012 	{int(X9)*1R}
R14 	N019 	N020 	{int(X10)*1R}
R15 	N019 	0 		{int(X11)*1R}
R16 	N006 	N007 	{int(X12)*1R}
R17 	N022 	0 		{int(X13)*1R}
R18 	N009 	N006 	{int(X14)*1R}
R28 	V_grid 	N004 	{int(X15)*1R}
R29 	N015 	V_grid 	{int(X16)*1R}
R32 	N016 	N015 	{int(X17)*1R}
R33 	N005 	N004 	{int(X18)*1R}


*LOAD RESISTOR
Rload 	0 		out 	8

*CAPACITORS
C1 		N010 	N009 	{int(X19)*1u}
C2 		N017 	N019 	{int(X20)*1n}
C3 		N022 	0 		{int(X21)*1u}
C5 		N015 	N008 	{int(X22)*1u}
C6 		N004 	N003 	{int(X23)*1u}

*BIPOLARS
Q1 	N013 N021 N023 	0 		BC847C
Q4 	N021 N023 0 	0 		BC847C

*OUTPUT TRANSFORMER
XU1 N001 N002 V_PP 	N014 	N018 out NC_01 0 PAT4002

*VALVES
XU2 N001 N002 N005 	0 		EL84
XU3 N018 N014 N016 	0 		EL84
XU6 N008 N011 N013 	12AU7
XU7 N003 N012 N013 	12AU7
XU8 V_PP N007 N009 	12AU7
XU9 N006 N020 N022 	12AU7

*SOURCES
V2 V_PP 0 {int(X24)}
V6 V_grid 0 {int(X25)}
B1 V_in 0 V=v(amp)*sin(2*pi*1000*time)
B2 amp 0 V={10m*ceil(time*100)-10m}
B3 tref 0 V={1*time}

*COMMANDS
.tran 0 1.01 0 10u
.probe v(out)
.MEAS TRAN MIN0 MIN V(out) FROM=0m TO=10m
.MEAS TRAN MAX0 MAX V(out) FROM=0m TO=10m
.MEAS TRAN MIN1 MIN V(out) FROM=10m TO=20m
.MEAS TRAN MAX1 MAX V(out) FROM=10m TO=20m
.MEAS TRAN MIN2 MIN V(out) FROM=20m TO=30m
.MEAS TRAN MAX2 MAX V(out) FROM=20m TO=30m
.MEAS TRAN MIN3 MIN V(out) FROM=30m TO=40m
.MEAS TRAN MAX3 MAX V(out) FROM=30m TO=40m
.MEAS TRAN MIN4 MIN V(out) FROM=40m TO=50m
.MEAS TRAN MAX4 MAX V(out) FROM=40m TO=50m
.MEAS TRAN MIN5 MIN V(out) FROM=50m TO=60m
.MEAS TRAN MAX5 MAX V(out) FROM=50m TO=60m
.MEAS TRAN MIN6 MIN V(out) FROM=60m TO=70m
.MEAS TRAN MAX6 MAX V(out) FROM=60m TO=70m
.MEAS TRAN MIN7 MIN V(out) FROM=70m TO=80m
.MEAS TRAN MAX7 MAX V(out) FROM=70m TO=80m
.MEAS TRAN MIN8 MIN V(out) FROM=80m TO=90m
.MEAS TRAN MAX8 MAX V(out) FROM=80m TO=90m
.MEAS TRAN MIN9 MIN V(out) FROM=90m TO=100m
.MEAS TRAN MAX9 MAX V(out) FROM=90m TO=100m
.MEAS TRAN MIN10 MIN V(out) FROM=100m TO=110m
.MEAS TRAN MAX10 MAX V(out) FROM=100m TO=110m
.MEAS TRAN MIN11 MIN V(out) FROM=110m TO=120m
.MEAS TRAN MAX11 MAX V(out) FROM=110m TO=120m
.MEAS TRAN MIN12 MIN V(out) FROM=120m TO=130m
.MEAS TRAN MAX12 MAX V(out) FROM=120m TO=130m
.MEAS TRAN MIN13 MIN V(out) FROM=130m TO=140m
.MEAS TRAN MAX13 MAX V(out) FROM=130m TO=140m
.MEAS TRAN MIN14 MIN V(out) FROM=140m TO=150m
.MEAS TRAN MAX14 MAX V(out) FROM=140m TO=150m
.MEAS TRAN MIN15 MIN V(out) FROM=150m TO=160m
.MEAS TRAN MAX15 MAX V(out) FROM=150m TO=160m
.MEAS TRAN MIN16 MIN V(out) FROM=160m TO=170m
.MEAS TRAN MAX16 MAX V(out) FROM=160m TO=170m
.MEAS TRAN MIN17 MIN V(out) FROM=170m TO=180m
.MEAS TRAN MAX17 MAX V(out) FROM=170m TO=180m
.MEAS TRAN MIN18 MIN V(out) FROM=180m TO=190m
.MEAS TRAN MAX18 MAX V(out) FROM=180m TO=190m
.MEAS TRAN MIN19 MIN V(out) FROM=190m TO=200m
.MEAS TRAN MAX19 MAX V(out) FROM=190m TO=200m
.MEAS TRAN MIN20 MIN V(out) FROM=200m TO=210m
.MEAS TRAN MAX20 MAX V(out) FROM=200m TO=210m
.MEAS TRAN MIN21 MIN V(out) FROM=210m TO=220m
.MEAS TRAN MAX21 MAX V(out) FROM=210m TO=220m
.MEAS TRAN MIN22 MIN V(out) FROM=220m TO=230m
.MEAS TRAN MAX22 MAX V(out) FROM=220m TO=230m
.MEAS TRAN MIN23 MIN V(out) FROM=230m TO=240m
.MEAS TRAN MAX23 MAX V(out) FROM=230m TO=240m
.MEAS TRAN MIN24 MIN V(out) FROM=240m TO=250m
.MEAS TRAN MAX24 MAX V(out) FROM=240m TO=250m
.MEAS TRAN MIN25 MIN V(out) FROM=250m TO=260m
.MEAS TRAN MAX25 MAX V(out) FROM=250m TO=260m
.MEAS TRAN MIN26 MIN V(out) FROM=260m TO=270m
.MEAS TRAN MAX26 MAX V(out) FROM=260m TO=270m
.MEAS TRAN MIN27 MIN V(out) FROM=270m TO=280m
.MEAS TRAN MAX27 MAX V(out) FROM=270m TO=280m
.MEAS TRAN MIN28 MIN V(out) FROM=280m TO=290m
.MEAS TRAN MAX28 MAX V(out) FROM=280m TO=290m
.MEAS TRAN MIN29 MIN V(out) FROM=290m TO=300m
.MEAS TRAN MAX29 MAX V(out) FROM=290m TO=300m
.MEAS TRAN MIN30 MIN V(out) FROM=300m TO=310m
.MEAS TRAN MAX30 MAX V(out) FROM=300m TO=310m
.MEAS TRAN MIN31 MIN V(out) FROM=310m TO=320m
.MEAS TRAN MAX31 MAX V(out) FROM=310m TO=320m
.MEAS TRAN MIN32 MIN V(out) FROM=320m TO=330m
.MEAS TRAN MAX32 MAX V(out) FROM=320m TO=330m
.MEAS TRAN MIN33 MIN V(out) FROM=330m TO=340m
.MEAS TRAN MAX33 MAX V(out) FROM=330m TO=340m
.MEAS TRAN MIN34 MIN V(out) FROM=340m TO=350m
.MEAS TRAN MAX34 MAX V(out) FROM=340m TO=350m
.MEAS TRAN MIN35 MIN V(out) FROM=350m TO=360m
.MEAS TRAN MAX35 MAX V(out) FROM=350m TO=360m
.MEAS TRAN MIN36 MIN V(out) FROM=360m TO=370m
.MEAS TRAN MAX36 MAX V(out) FROM=360m TO=370m
.MEAS TRAN MIN37 MIN V(out) FROM=370m TO=380m
.MEAS TRAN MAX37 MAX V(out) FROM=370m TO=380m
.MEAS TRAN MIN38 MIN V(out) FROM=380m TO=390m
.MEAS TRAN MAX38 MAX V(out) FROM=380m TO=390m
.MEAS TRAN MIN39 MIN V(out) FROM=390m TO=400m
.MEAS TRAN MAX39 MAX V(out) FROM=390m TO=400m
.MEAS TRAN MIN40 MIN V(out) FROM=400m TO=410m
.MEAS TRAN MAX40 MAX V(out) FROM=400m TO=410m
.MEAS TRAN MIN41 MIN V(out) FROM=410m TO=420m
.MEAS TRAN MAX41 MAX V(out) FROM=410m TO=420m
.MEAS TRAN MIN42 MIN V(out) FROM=420m TO=430m
.MEAS TRAN MAX42 MAX V(out) FROM=420m TO=430m
.MEAS TRAN MIN43 MIN V(out) FROM=430m TO=440m
.MEAS TRAN MAX43 MAX V(out) FROM=430m TO=440m
.MEAS TRAN MIN44 MIN V(out) FROM=440m TO=450m
.MEAS TRAN MAX44 MAX V(out) FROM=440m TO=450m
.MEAS TRAN MIN45 MIN V(out) FROM=450m TO=460m
.MEAS TRAN MAX45 MAX V(out) FROM=450m TO=460m
.MEAS TRAN MIN46 MIN V(out) FROM=460m TO=470m
.MEAS TRAN MAX46 MAX V(out) FROM=460m TO=470m
.MEAS TRAN MIN47 MIN V(out) FROM=470m TO=480m
.MEAS TRAN MAX47 MAX V(out) FROM=470m TO=480m
.MEAS TRAN MIN48 MIN V(out) FROM=480m TO=490m
.MEAS TRAN MAX48 MAX V(out) FROM=480m TO=490m
.MEAS TRAN MIN49 MIN V(out) FROM=490m TO=500m
.MEAS TRAN MAX49 MAX V(out) FROM=490m TO=500m
.MEAS TRAN MIN50 MIN V(out) FROM=500m TO=510m
.MEAS TRAN MAX50 MAX V(out) FROM=500m TO=510m
.MEAS TRAN MIN51 MIN V(out) FROM=510m TO=520m
.MEAS TRAN MAX51 MAX V(out) FROM=510m TO=520m
.MEAS TRAN MIN52 MIN V(out) FROM=520m TO=530m
.MEAS TRAN MAX52 MAX V(out) FROM=520m TO=530m
.MEAS TRAN MIN53 MIN V(out) FROM=530m TO=540m
.MEAS TRAN MAX53 MAX V(out) FROM=530m TO=540m
.MEAS TRAN MIN54 MIN V(out) FROM=540m TO=550m
.MEAS TRAN MAX54 MAX V(out) FROM=540m TO=550m
.MEAS TRAN MIN55 MIN V(out) FROM=550m TO=560m
.MEAS TRAN MAX55 MAX V(out) FROM=550m TO=560m
.MEAS TRAN MIN56 MIN V(out) FROM=560m TO=570m
.MEAS TRAN MAX56 MAX V(out) FROM=560m TO=570m
.MEAS TRAN MIN57 MIN V(out) FROM=570m TO=580m
.MEAS TRAN MAX57 MAX V(out) FROM=570m TO=580m
.MEAS TRAN MIN58 MIN V(out) FROM=580m TO=590m
.MEAS TRAN MAX58 MAX V(out) FROM=580m TO=590m
.MEAS TRAN MIN59 MIN V(out) FROM=590m TO=600m
.MEAS TRAN MAX59 MAX V(out) FROM=590m TO=600m
.MEAS TRAN MIN60 MIN V(out) FROM=600m TO=610m
.MEAS TRAN MAX60 MAX V(out) FROM=600m TO=610m
.MEAS TRAN MIN61 MIN V(out) FROM=610m TO=620m
.MEAS TRAN MAX61 MAX V(out) FROM=610m TO=620m
.MEAS TRAN MIN62 MIN V(out) FROM=620m TO=630m
.MEAS TRAN MAX62 MAX V(out) FROM=620m TO=630m
.MEAS TRAN MIN63 MIN V(out) FROM=630m TO=640m
.MEAS TRAN MAX63 MAX V(out) FROM=630m TO=640m
.MEAS TRAN MIN64 MIN V(out) FROM=640m TO=650m
.MEAS TRAN MAX64 MAX V(out) FROM=640m TO=650m
.MEAS TRAN MIN65 MIN V(out) FROM=650m TO=660m
.MEAS TRAN MAX65 MAX V(out) FROM=650m TO=660m
.MEAS TRAN MIN66 MIN V(out) FROM=660m TO=670m
.MEAS TRAN MAX66 MAX V(out) FROM=660m TO=670m
.MEAS TRAN MIN67 MIN V(out) FROM=670m TO=680m
.MEAS TRAN MAX67 MAX V(out) FROM=670m TO=680m
.MEAS TRAN MIN68 MIN V(out) FROM=680m TO=690m
.MEAS TRAN MAX68 MAX V(out) FROM=680m TO=690m
.MEAS TRAN MIN69 MIN V(out) FROM=690m TO=700m
.MEAS TRAN MAX69 MAX V(out) FROM=690m TO=700m
.MEAS TRAN MIN70 MIN V(out) FROM=700m TO=710m
.MEAS TRAN MAX70 MAX V(out) FROM=700m TO=710m
.MEAS TRAN MIN71 MIN V(out) FROM=710m TO=720m
.MEAS TRAN MAX71 MAX V(out) FROM=710m TO=720m
.MEAS TRAN MIN72 MIN V(out) FROM=720m TO=730m
.MEAS TRAN MAX72 MAX V(out) FROM=720m TO=730m
.MEAS TRAN MIN73 MIN V(out) FROM=730m TO=740m
.MEAS TRAN MAX73 MAX V(out) FROM=730m TO=740m
.MEAS TRAN MIN74 MIN V(out) FROM=740m TO=750m
.MEAS TRAN MAX74 MAX V(out) FROM=740m TO=750m
.MEAS TRAN MIN75 MIN V(out) FROM=750m TO=760m
.MEAS TRAN MAX75 MAX V(out) FROM=750m TO=760m
.MEAS TRAN MIN76 MIN V(out) FROM=760m TO=770m
.MEAS TRAN MAX76 MAX V(out) FROM=760m TO=770m
.MEAS TRAN MIN77 MIN V(out) FROM=770m TO=780m
.MEAS TRAN MAX77 MAX V(out) FROM=770m TO=780m
.MEAS TRAN MIN78 MIN V(out) FROM=780m TO=790m
.MEAS TRAN MAX78 MAX V(out) FROM=780m TO=790m
.MEAS TRAN MIN79 MIN V(out) FROM=790m TO=800m
.MEAS TRAN MAX79 MAX V(out) FROM=790m TO=800m
.MEAS TRAN MIN80 MIN V(out) FROM=800m TO=810m
.MEAS TRAN MAX80 MAX V(out) FROM=800m TO=810m
.MEAS TRAN MIN81 MIN V(out) FROM=810m TO=820m
.MEAS TRAN MAX81 MAX V(out) FROM=810m TO=820m
.MEAS TRAN MIN82 MIN V(out) FROM=820m TO=830m
.MEAS TRAN MAX82 MAX V(out) FROM=820m TO=830m
.MEAS TRAN MIN83 MIN V(out) FROM=830m TO=840m
.MEAS TRAN MAX83 MAX V(out) FROM=830m TO=840m
.MEAS TRAN MIN84 MIN V(out) FROM=840m TO=850m
.MEAS TRAN MAX84 MAX V(out) FROM=840m TO=850m
.MEAS TRAN MIN85 MIN V(out) FROM=850m TO=860m
.MEAS TRAN MAX85 MAX V(out) FROM=850m TO=860m
.MEAS TRAN MIN86 MIN V(out) FROM=860m TO=870m
.MEAS TRAN MAX86 MAX V(out) FROM=860m TO=870m
.MEAS TRAN MIN87 MIN V(out) FROM=870m TO=880m
.MEAS TRAN MAX87 MAX V(out) FROM=870m TO=880m
.MEAS TRAN MIN88 MIN V(out) FROM=880m TO=890m
.MEAS TRAN MAX88 MAX V(out) FROM=880m TO=890m
.MEAS TRAN MIN89 MIN V(out) FROM=890m TO=900m
.MEAS TRAN MAX89 MAX V(out) FROM=890m TO=900m
.MEAS TRAN MIN90 MIN V(out) FROM=900m TO=910m
.MEAS TRAN MAX90 MAX V(out) FROM=900m TO=910m
.MEAS TRAN MIN91 MIN V(out) FROM=910m TO=920m
.MEAS TRAN MAX91 MAX V(out) FROM=910m TO=920m
.MEAS TRAN MIN92 MIN V(out) FROM=920m TO=930m
.MEAS TRAN MAX92 MAX V(out) FROM=920m TO=930m
.MEAS TRAN MIN93 MIN V(out) FROM=930m TO=940m
.MEAS TRAN MAX93 MAX V(out) FROM=930m TO=940m
.MEAS TRAN MIN94 MIN V(out) FROM=940m TO=950m
.MEAS TRAN MAX94 MAX V(out) FROM=940m TO=950m
.MEAS TRAN MIN95 MIN V(out) FROM=950m TO=960m
.MEAS TRAN MAX95 MAX V(out) FROM=950m TO=960m
.MEAS TRAN MIN96 MIN V(out) FROM=960m TO=970m
.MEAS TRAN MAX96 MAX V(out) FROM=960m TO=970m
.MEAS TRAN MIN97 MIN V(out) FROM=970m TO=980m
.MEAS TRAN MAX97 MAX V(out) FROM=970m TO=980m
.MEAS TRAN MIN98 MIN V(out) FROM=980m TO=990m
.MEAS TRAN MAX98 MAX V(out) FROM=980m TO=990m
.MEAS TRAN MIN99 MIN V(out) FROM=990m TO=1000m
.MEAS TRAN MAX99 MAX V(out) FROM=990m TO=1000m
.MEAS TRAN MIN100 MIN V(out) FROM=1000m TO=1010m
.MEAS TRAN MAX100 MAX V(out) FROM=1000m TO=1010m


*INCLUDES
.include ./param.txt
.model NPN NPN
.model PNP PNP
.lib C:\Users\Colombari\Documents\LTspiceXVII\lib\cmp\standard.bjt
.lib trafos.lib
.lib tube.lib
.lib tubes.lib
.backanno
.end
